`include "core.sv"

module test();


endmodule