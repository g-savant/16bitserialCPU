module instr_shift_register(

);

endmodule


module instruction_decode(
  input logic[15:0] instruction,
  output signals_t signals
);

  always_comb begin
    signals.opcode = 
  end

endmodule