// `default_nettype none

// module Counter(

// );

// endmodule