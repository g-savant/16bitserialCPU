module test();





endmodule